// $Id: $
// File name:   tb_horizontal_gradient.sv
// Created:     4/22/2016
// Author:
// Lab Section: 337-01
// Version:     1.0  Initial Design Entry
// Description: tb for horizontal_gradient.sv
`timescale 1ns / 100ps

module tb_horizontal_gradient ();
  
  
