module check_edge(

input wire [7:0] G,
output reg calculation_done,
output reg [7:0] edge

);

  //check edge here return 0 or 255 depending on the value of G 
  
  
  
  
endmodule
