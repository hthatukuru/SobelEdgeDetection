module check_edge(

input wire [7:0] G,
output reg calculation_done,
output reg [7:0] edge


);
