// $Id: $
// File name:   tb_vertical_gradient.sv
// Created:     4/22/2016
// Author:   
// Lab Section: 337-01
// Version:     1.0  Initial Design Entry
// Description: tb for vertical_gradient.sv
`timescale 1ns / 100ps
