module ahb_slave(
output reg start,
output reg [11:0] width, length,
output reg [7:0] initial_addr_r, initial_addr_w,
);





endmodule
